`timescale 1ns/10ps
//////////////////////////////////////////////////////////////////////////////////
// Company:         Tel Aviv University
// Engineer:        
// 
// Create Date:     05/05/2019 02:59:38 AM
// Design Name:     EE3 lab1
// Module Name:     Ctl_tb
// Project Name:    Electrical Lab 3, FPGA Experiment #1
// Target Devices:  Xilinx BASYS3 Board, FPGA model XC7A35T-lcpg236C
// Tool versions:   Vivado 2016.4
// Description:     test bennch for the control.
// Dependencies:    None
//
// Revision: 		3.0
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module Ctl_tb();

    reg clk, reset, trig, split, correct;
    wire init_regs, count_enabled;
    //integer ai,cii;
    
    // Instantiate the UUT (Unit Under Test)
    Ctl uut (clk, reset, trig, split, init_regs, count_enabled);
    // FILL HERE
    initial begin
        correct = 1;
        clk = 0; 
        reset = 1; 
        trig = 0;
        split = 0;
        #10
        reset = 0; 
        correct = correct & init_regs & ~count_enabled;
        #20
        trig = 1;
        #10
        trig = 0;
        #10
        correct = correct & (~init_regs) & (count_enabled);
        trig = 1;
        #10
        trig = 0;
        #10
        correct = correct & (~init_regs) & (~count_enabled);
        trig = 1;
        #20
        trig = 0;
        #10
        split = 1;
        #10
        split = 0;
        #10
        correct = correct & (init_regs) & (~count_enabled);
        #10
        if (correct)
            $display("Test Passed - %m");
        else
            $display("Test Failed - %m");
        $finish;
    end
    
    always #5 clk = ~clk;
    
endmodule
